* # FILE NAME: /NFS/STAK/STUDENTS/B/BRANAUGJ/CADENCE/SIMULATION/LAB6_CLA/       
* HSPICES/SCHEMATIC/NETLIST/LAB6_CLA.C.RAW
* NETLIST OUTPUT FOR HSPICES.
* GENERATED ON FEB 28 15:26:50 2014
   
* GLOBAL NET DEFINITIONS
.GLOBAL VDD! 
* FILE NAME: ECE471_LIB_LAB6_CLA_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: LAB6_CLA.
* GENERATED FOR: HSPICES.
* GENERATED ON FEB 28 15:26:51 2014.
   
XI4 A0 B0 C0 NET28 NET50 NET46 S0 SUB1 
XI3 A1 B1 NET55 NET35 NET49 NET45 S1 SUB1 
XI2 A2 B2 NET36 NET42 NET41 NET40 S2 SUB1 
XI1 A3 B3 NET15 NET21 NET20 NET19 S3 SUB1 
XI0 C0 NET55 NET36 NET15 C4 NET50 NET49 NET41 NET20 NET46 NET45 NET40 NET19 
+SUB2 
   
   
   
   
* FILE NAME: ECE471_LIB_LAB6_FULL_ADDER_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: LAB6_FULL_ADDER.
* GENERATED FOR: HSPICES.
* GENERATED ON FEB 28 15:26:51 2014.
   
* TERMINAL MAPPING: AI = AI
*                   BI = BI
*                   CI = CI
*                   CO = CO
*                   GI = GI
*                   PI = PI
*                   SI = SI
.SUBCKT SUB1 AI BI CI CO GI PI SI 
XI5 GI NET09 CO OR2_1 
XI3 AI BI PI LAB6_XOR_G1 
XI2 CI AI NET018 LAB6_XOR_G1 
XI1 NET018 BI SI LAB6_XOR_G1 
XI4 PI CI NET09 AND2_2 
XI0 AI BI GI AND2_2 
   
   
* FILE NAME: NCSU_DIGITAL_PARTS_AND2_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: AND2.
* GENERATED FOR: HSPICES.
* GENERATED ON FEB 28 15:26:51 2014.
   
* TERMINAL MAPPING: A = A
*                   B = B
*                   Y = Y
.SUBCKT AND2_2 A B Y 
M5 Y NET29 VDD! VDD!  TSMC25DP  L=(240E-9) W=(720E-9) AD=+4.32000000E-13 
+AS=+4.32000000E-13 PD=+2.64000000E-06 PS=+2.64000000E-06 OFF 
M3 NET29 B VDD! VDD!  TSMC25DP  L=(240E-9) W=(720E-9) AD=+4.32000000E-13 
+AS=+4.32000000E-13 PD=+2.64000000E-06 PS=+2.64000000E-06 OFF 
M2 NET29 A VDD! VDD!  TSMC25DP  L=(240E-9) W=(720E-9) AD=+4.32000000E-13 
+AS=+4.32000000E-13 PD=+2.64000000E-06 PS=+2.64000000E-06 OFF 
M4 Y NET29 0 0  TSMC25DN  L=(240E-9) W=(360E-9) AD=+2.16000000E-13 
+AS=+2.16000000E-13 PD=+1.92000000E-06 PS=+1.92000000E-06 OFF 
M1 NET29 A NET11 0  TSMC25DN  L=(240E-9) W=(360E-9) AD=+2.16000000E-13 
+AS=+2.16000000E-13 PD=+1.92000000E-06 PS=+1.92000000E-06 OFF 
M0 NET11 B 0 0  TSMC25DN  L=(240E-9) W=(360E-9) AD=+2.16000000E-13 
+AS=+2.16000000E-13 PD=+1.92000000E-06 PS=+1.92000000E-06 OFF 
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS AND2_2 
* FILE NAME: NCSU_DIGITAL_PARTS_OR2_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: OR2.
* GENERATED FOR: HSPICES.
* GENERATED ON FEB 28 15:26:50 2014.
   
* TERMINAL MAPPING: A = A
*                   B = B
*                   Y = Y
.SUBCKT OR2_1 A B Y 
M5 Y NET21 VDD! VDD!  TSMC25DP  L=(240E-9) W=(1.44E-6) AD=+8.64000000E-13 
+AS=+8.64000000E-13 PD=+4.08000000E-06 PS=+4.08000000E-06 OFF 
M3 NET11 A VDD! VDD!  TSMC25DP  L=(240E-9) W=(1.44E-6) AD=+8.64000000E-13 
+AS=+8.64000000E-13 PD=+4.08000000E-06 PS=+4.08000000E-06 OFF 
M2 NET21 B NET11 VDD!  TSMC25DP  L=(240E-9) W=(1.44E-6) AD=+8.64000000E-13 
+AS=+8.64000000E-13 PD=+4.08000000E-06 PS=+4.08000000E-06 OFF 
M4 Y NET21 0 0  TSMC25DN  L=(240E-9) W=(360E-9) AD=+2.16000000E-13 
+AS=+2.16000000E-13 PD=+1.92000000E-06 PS=+1.92000000E-06 OFF 
M1 NET21 B 0 0  TSMC25DN  L=(240E-9) W=(360E-9) AD=+2.16000000E-13 
+AS=+2.16000000E-13 PD=+1.92000000E-06 PS=+1.92000000E-06 OFF 
M0 NET21 A 0 0  TSMC25DN  L=(240E-9) W=(360E-9) AD=+2.16000000E-13 
+AS=+2.16000000E-13 PD=+1.92000000E-06 PS=+1.92000000E-06 OFF 
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS OR2_1 
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SUB1 
* FILE NAME: ECE471_LIB_LAB6_XOR_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: LAB6_XOR.
* GENERATED FOR: HSPICES.
* GENERATED ON FEB 28 15:26:51 2014.
   
* TERMINAL MAPPING: A = A
*                   B = B
*                   Y = Y
.SUBCKT LAB6_XOR_G1 A B Y 
MN5 1 B 0 0  TSMC25DN  L=240E-9 W=360E-9 AD=216E-15 AS=216E-15 PD=1.92E-6 
+PS=1.92E-6 M=1 
MN4 2 A 0 0  TSMC25DN  L=240E-9 W=360E-9 AD=216E-15 AS=216E-15 PD=1.92E-6 
+PS=1.92E-6 M=1 
MN3 NET12 1 0 0  TSMC25DN  L=240E-9 W=720E-9 AD=432E-15 AS=432E-15 PD=2.64E-6 
+PS=2.64E-6 M=1 
MN2 NET16 B 0 0  TSMC25DN  L=240E-9 W=720E-9 AD=432E-15 AS=432E-15 PD=2.64E-6 
+PS=2.64E-6 M=1 
MN1 Y A NET16 0  TSMC25DN  L=240E-9 W=720E-9 AD=432E-15 AS=432E-15 PD=2.64E-6 
+PS=2.64E-6 M=1 
MN0 Y 2 NET12 0  TSMC25DN  L=240E-9 W=720E-9 AD=432E-15 AS=432E-15 PD=2.64E-6 
+PS=2.64E-6 M=1 
MP5 1 B VDD! VDD!  TSMC25DP  L=240E-9 W=720E-9 AD=432E-15 AS=432E-15 
+PD=2.64E-6 PS=2.64E-6 M=1 
MP4 2 A VDD! VDD!  TSMC25DP  L=240E-9 W=720E-9 AD=432E-15 AS=432E-15 
+PD=2.64E-6 PS=2.64E-6 M=1 
MP3 Y 1 NET47 VDD!  TSMC25DP  L=240E-9 W=1.44E-6 AD=864E-15 AS=864E-15 
+PD=4.08E-6 PS=4.08E-6 M=1 
MP2 NET47 B VDD! VDD!  TSMC25DP  L=240E-9 W=1.44E-6 AD=864E-15 AS=864E-15 
+PD=4.08E-6 PS=4.08E-6 M=1 
MP1 Y 2 NET47 VDD!  TSMC25DP  L=240E-9 W=1.44E-6 AD=864E-15 AS=864E-15 
+PD=4.08E-6 PS=4.08E-6 M=1 
MP0 NET47 A VDD! VDD!  TSMC25DP  L=240E-9 W=1.44E-6 AD=864E-15 AS=864E-15 
+PD=4.08E-6 PS=4.08E-6 M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS LAB6_XOR_G1 
* FILE NAME: ECE471_LIB_LAB6_CARRY_BLOCK_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: LAB6_CARRY_BLOCK.
* GENERATED FOR: HSPICES.
* GENERATED ON FEB 28 15:26:51 2014.
   
* TERMINAL MAPPING: C0 = C0
*                   C1 = C1
*                   C2 = C2
*                   C3 = C3
*                   C4 = C4
*                   G0 = G0
*                   G1 = G1
*                   G2 = G2
*                   G3 = G3
*                   P0 = P0
*                   P1 = P1
*                   P2 = P2
*                   P3 = P3
.SUBCKT SUB2 C0 C1 C2 C3 C4 G0 G1 G2 G3 P0 P1 P2 P3 
XI16 G0 NET064 NET034 OR2_1 
XI14 G2 NET070 NET040 OR2_1 
XI15 G1 NET067 NET037 OR2_1 
XI10 G0 NET079 NET049 OR2_1 
XI11 G1 NET076 NET046 OR2_1 
XI8 G0 NET082 NET052 OR2_1 
XI5 G3 NET26 C4 OR2_1 
XI4 G2 NET29 C3 OR2_1 
XI1 G0 NET35 C1 OR2_1 
XI3 G1 NET32 C2 OR2_1 
XI19 C0 P0 NET064 AND2_2 
XI18 NET034 P1 NET067 AND2_2 
XI17 NET037 P2 NET070 AND2_2 
XI12 C0 P0 NET079 AND2_2 
XI13 NET049 P1 NET076 AND2_2 
XI7 NET040 P3 NET26 AND2_2 
XI6 NET046 P2 NET29 AND2_2 
XI2 NET052 P1 NET32 AND2_2 
XI0 C0 P0 NET35 AND2_2 
XI9 C0 P0 NET082 AND2_2 
   
   
* FILE NAME: NCSU_DIGITAL_PARTS_OR2_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: OR2.
* GENERATED FOR: HSPICES.
* GENERATED ON FEB 28 15:26:50 2014.
   
* TERMINAL MAPPING: A = A
*                   B = B
*                   Y = Y
.SUBCKT OR2_1 A B Y 
M5 Y NET21 VDD! VDD!  TSMC25DP  L=(240E-9) W=(2.88E-6) AD=+1.72800000E-12 
+AS=+1.72800000E-12 PD=+6.96000000E-06 PS=+6.96000000E-06 OFF 
M3 NET11 A VDD! VDD!  TSMC25DP  L=(240E-9) W=(2.88E-6) AD=+1.72800000E-12 
+AS=+1.72800000E-12 PD=+6.96000000E-06 PS=+6.96000000E-06 OFF 
M2 NET21 B NET11 VDD!  TSMC25DP  L=(240E-9) W=(2.88E-6) AD=+1.72800000E-12 
+AS=+1.72800000E-12 PD=+6.96000000E-06 PS=+6.96000000E-06 OFF 
M4 Y NET21 0 0  TSMC25DN  L=(240E-9) W=(1.44E-6) AD=+8.64000000E-13 
+AS=+8.64000000E-13 PD=+4.08000000E-06 PS=+4.08000000E-06 OFF 
M1 NET21 B 0 0  TSMC25DN  L=(240E-9) W=(1.44E-6) AD=+8.64000000E-13 
+AS=+8.64000000E-13 PD=+4.08000000E-06 PS=+4.08000000E-06 OFF 
M0 NET21 A 0 0  TSMC25DN  L=(240E-9) W=(1.44E-6) AD=+8.64000000E-13 
+AS=+8.64000000E-13 PD=+4.08000000E-06 PS=+4.08000000E-06 OFF 
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS OR2_1 
* FILE NAME: NCSU_DIGITAL_PARTS_AND2_CMOS_SCH.S.
* SUBCIRCUIT FOR CELL: AND2.
* GENERATED FOR: HSPICES.
* GENERATED ON FEB 28 15:26:51 2014.
   
* TERMINAL MAPPING: A = A
*                   B = B
*                   Y = Y
.SUBCKT AND2_2 A B Y 
M5 Y NET29 VDD! VDD!  TSMC25DP  L=(240E-9) W=(2.88E-6) AD=+1.72800000E-12 
+AS=+1.72800000E-12 PD=+6.96000000E-06 PS=+6.96000000E-06 OFF 
M3 NET29 B VDD! VDD!  TSMC25DP  L=(240E-9) W=(2.88E-6) AD=+1.72800000E-12 
+AS=+1.72800000E-12 PD=+6.96000000E-06 PS=+6.96000000E-06 OFF 
M2 NET29 A VDD! VDD!  TSMC25DP  L=(240E-9) W=(2.88E-6) AD=+1.72800000E-12 
+AS=+1.72800000E-12 PD=+6.96000000E-06 PS=+6.96000000E-06 OFF 
M4 Y NET29 0 0  TSMC25DN  L=(240E-9) W=(1.44E-6) AD=+8.64000000E-13 
+AS=+8.64000000E-13 PD=+4.08000000E-06 PS=+4.08000000E-06 OFF 
M1 NET29 A NET11 0  TSMC25DN  L=(240E-9) W=(1.44E-6) AD=+8.64000000E-13 
+AS=+8.64000000E-13 PD=+4.08000000E-06 PS=+4.08000000E-06 OFF 
M0 NET11 B 0 0  TSMC25DN  L=(240E-9) W=(1.44E-6) AD=+8.64000000E-13 
+AS=+8.64000000E-13 PD=+4.08000000E-06 PS=+4.08000000E-06 OFF 
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS AND2_2 
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SUB2 
