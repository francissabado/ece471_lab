* # FILE NAME: /NFS/STAK/STUDENTS/B/BRANAUGJ/CADENCE/SIMULATION/LAB3_CKT/       
* HSPICES/SCHEMATIC/NETLIST/LAB3_CKT.C.RAW
* NETLIST OUTPUT FOR HSPICES.
* GENERATED ON JAN 31 15:30:11 2014
   
* GLOBAL NET DEFINITIONS
.GLOBAL VDD! GND! 
* FILE NAME: ECE471_LIB_LAB3_CKT_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: LAB3_CKT.
* GENERATED FOR: HSPICES.
* GENERATED ON JAN 31 15:30:11 2014.
   
R2 NET4 NET07  6.53 M=1.0 
R3 NET03 NET05  6.53 M=1.0 
R0 NET07 NET03  6.53 M=1.0 
C2 NET05 GND!  8.41E-15 M=1.0 
C3 NET4 GND!  8.41E-15 M=1.0 
C0 NET07 GND!  16.83E-15 M=1.0 
C1 NET03 GND!  16.83E-15 M=1.0 
XI2 VIN NET4 INVERTER_G1 
XI3 NET05 VOUT INVERTER_G1 
   
   
   
   
* FILE NAME: ECE471_LIB_INVERTER_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: INVERTER.
* GENERATED FOR: HSPICES.
* GENERATED ON JAN 31 15:30:11 2014.
   
* TERMINAL MAPPING: INPUT = INPUT
*                   OUTPUT = OUTPUT
.SUBCKT INVERTER_G1 INPUT OUTPUT 
MP0 OUTPUT INPUT VDD! VDD!  TSMC25DP  L=240E-9 W=960E-9 AD=576E-15 AS=576E-15 
+PD=3.12E-6 PS=3.12E-6 M=1 
MN0 OUTPUT INPUT 0 0  TSMC25DN  L=240E-9 W=480E-9 AD=288E-15 AS=288E-15 
+PD=2.16E-6 PS=2.16E-6 M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INVERTER_G1 
